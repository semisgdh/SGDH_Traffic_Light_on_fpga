// common_defines.vh
`define TIMER_BIT_WIDTH 32

// timescale definition
`timescale 1ns/1ps